--Christos Gkoumas, p3160026
--Spyridon Pagkalos, p3150133

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--PACKAGE DECLARATION FOR ALL THE REQUIRED SUBCIRCUITS
PACKAGE subcircuits IS
	--COMPONENT DECLARATION FOR 16-BIT AND
	COMPONENT GATE_AND PORT (A, B: IN STD_LOGIC_VECTOR (15 DOWNTO 0); O: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
	END COMPONENT;
	--COMPONENT DECLARATION FOR 16-BIT OR
	COMPONENT GATE_OR PORT (A, B: IN STD_LOGIC_VECTOR (15 DOWNTO 0); O: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
	END COMPONENT;
	--COMPONENT DECLARATION FOR 16-BIT GEQ
	COMPONENT GATE_GEQ PORT (A: IN STD_LOGIC_VECTOR (15 DOWNTO 0); O: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
	END COMPONENT;
	--COMPONENT DECLARATION FOR 16-BIT NOT THAT IS ASKED IN THE PROJECT
	COMPONENT GATE_PR_NOT PORT (A: IN STD_LOGIC_VECTOR (15 DOWNTO 0); O:  OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
	END COMPONENT;
	--COMPONENT DECLARATION FOR 1-BIT AND
	COMPONENT GATE_AND_2 PORT (A, B: IN STD_LOGIC; O: OUT STD_LOGIC);
	END COMPONENT;
	--COMPONENT DECLARATION FOR 1-BIT OR WITH 3 INPUTS
	COMPONENT GATE_OR_3 PORT (A, B, C: IN STD_LOGIC; O: OUT STD_LOGIC);
	END COMPONENT;
	--COMPONENT DECLARATION FOR 1-BIT XOR
	COMPONENT GATE_XOR PORT (A, B: IN STD_LOGIC; O: OUT STD_LOGIC);
	END COMPONENT;
	--COMPONENT DECLARATION FOR 1-BIT XOR WITH 3 INPUTS
	COMPONENT GATE_XOR_3 PORT (A, B, C: IN STD_LOGIC; O: OUT STD_LOGIC);
	END COMPONENT;
	--COMPONENT DECLARATION FOR 1-BIT NOT
	COMPONENT GATE_NOT PORT (A: IN STD_LOGIC; O: OUT STD_LOGIC);
	END COMPONENT;
	--COMPONENT DECLARATION FOR 16-BIT NOT
	COMPONENT GATE_NOT_16 PORT (A: IN STD_LOGIC_VECTOR(15 DOWNTO 0); O: OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
	END COMPONENT;
	--COMPONENT DECLARATION FOR 1-BIT ADDER
	COMPONENT FULLADDER PORT(A, B, CIN: IN STD_LOGIC; O, COUT: OUT STD_LOGIC);
	END COMPONENT;
	--COMPONENT DECLARATION FOR 16-BIT ADDER
	COMPONENT FULLADDER_16 PORT(A, B: IN STD_LOGIC_VECTOR (15 DOWNTO 0); CIN: IN STD_LOGIC; O16: OUT STD_LOGIC_VECTOR (15 DOWNTO 0); V, COUT: OUT STD_LOGIC);
	END COMPONENT;
	--COMPONENT DECLARATION FOR 16-BIT SUBTRACTOR
	COMPONENT SUBTRACTOR_16 PORT(A, B: IN STD_LOGIC_VECTOR (15 DOWNTO 0); CIN: IN STD_LOGIC; O16: OUT STD_LOGIC_VECTOR (15 DOWNTO 0); V, COUT: OUT STD_LOGIC);
	END COMPONENT;
	--COMPONENT DECLARATION FOR COUNTER
	COMPONENT COUNTER PORT(CLEAR, CLOCK: IN STD_LOGIC; Q: BUFFER STD_LOGIC_VECTOR(1 DOWNTO 0));
	END COMPONENT;
	--COMPONENT DECLARATION FOR 16-BIT FLIP FLOP
	COMPONENT REG PORT (I: IN STD_LOGIC_VECTOR(15 DOWNTO 0); EN, CLOCK: IN STD_LOGIC; O: BUFFER STD_LOGIC_VECTOR(15 DOWNTO 0));
	END COMPONENT;
END PACKAGE;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--ENTITY DECLARATION FOR 16-BIT AND
ENTITY GATE_AND IS
	PORT (A, B: IN STD_LOGIC_VECTOR (15 DOWNTO 0); O: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END GATE_AND;

--ARCHITECTURE DECLARATION FOR 16-BIT AND
ARCHITECTURE Structural OF GATE_AND IS BEGIN
	O <= A AND B;
END Structural;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--ENTITY DECLARATION FOR 16-BIT OR
ENTITY GATE_OR IS
	PORT (A, B: IN STD_LOGIC_VECTOR (15 DOWNTO 0); O: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END GATE_OR;

--ARCHITECTURE DECLARATION FOR 16-BIT AND
ARCHITECTURE Structural OF GATE_OR IS BEGIN
	O <= A OR B;
END Structural;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--ENTITY DECLARATION FOR 16-BIT GEQ
ENTITY GATE_GEQ IS
	PORT (A: IN STD_LOGIC_VECTOR (15 DOWNTO 0); O: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END GATE_GEQ;

--ARCHITECTURE DECLARATION FOR 16-BIT AND
ARCHITECTURE Structural OF GATE_GEQ IS
SIGNAL TOUT: STD_LOGIC_VECTOR (15 DOWNTO 0);
BEGIN
	PROCESS(A)
	BEGIN
		IF (A(15)='0') THEN
			TOUT <= "1111111111111111";
		ELSE
			TOUT <= "0000000000000000";
		END IF;
		O <= TOUT;
	END PROCESS;
END Structural;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--ENTITY DECLARATION FOR 16-BIT NOT THAT IS ASKED IN THE PROJECT
ENTITY GATE_PR_NOT IS
	PORT (A: IN STD_LOGIC_VECTOR (15 DOWNTO 0); O: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END GATE_PR_NOT;

--ARCHITECTURE DECLARATION FOR 16-BIT NOT THAT IS ASKED IN THE PROJECT
ARCHITECTURE Structural OF GATE_PR_NOT IS
SIGNAL TOUT: STD_LOGIC_VECTOR (15 DOWNTO 0);
BEGIN
	PROCESS(A)
	BEGIN
		IF (A(0)= '1') THEN
			FOR I IN 1 TO 15 LOOP
				IF (A(I)/='0') THEN
					TOUT <= "0000000000000000";
					EXIT;
				END IF;
				TOUT <= "1111111111111111";
			END LOOP;
		ELSE
			TOUT <= "0000000000000000";
		END IF;
		O <= TOUT;
	END PROCESS;
END Structural;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--ENTITY DECLARATION FOR 1-BIT AND
ENTITY GATE_AND_2 IS
	PORT (A, B: IN STD_LOGIC; O: OUT STD_LOGIC);
END GATE_AND_2;

--ARCHITECTURE DECLARATION FOR 1-BIT AND
ARCHITECTURE Structural OF GATE_AND_2 IS 
BEGIN
	O <= A AND B;
END Structural;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--ENTITY DECLARATION FOR 1-BIT OR WITH 3 INPUTS
ENTITY GATE_OR_3 IS
	PORT (A, B, C: IN STD_LOGIC; O: OUT STD_LOGIC);
END GATE_OR_3;

--ARCHITECTURE DECLARATION FOR 1-BIT OR WITH 3 INPUTS
ARCHITECTURE Structural OF GATE_OR_3 IS
BEGIN
	O <= A OR B OR C;
END Structural;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--ENTITY DECLARATION FOR 1-BIT XOR
ENTITY GATE_XOR IS
	PORT (A, B: IN STD_LOGIC; O: OUT STD_LOGIC);
END GATE_XOR;

--ARCHITECTURE DECLARATION FOR 1-BIT XOR WITH 3 INPUTS
ARCHITECTURE Structural OF GATE_XOR IS BEGIN
	O <= A XOR B;
END Structural;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--ENTITY DECLARATION FOR 1-BIT XOR WITH 3 INPUTS
ENTITY GATE_XOR_3 IS
	PORT (A, B, C: IN STD_LOGIC; O: OUT STD_LOGIC);
END GATE_XOR_3;

--ARCHITECTURE DECLARATION FOR 1-BIT XOR WITH 3 INPUTS
ARCHITECTURE Structural OF GATE_XOR_3 IS BEGIN
	O <= A XOR B XOR C;
END Structural;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--ENTITY DECLARATION FOR 1-BIT NOT
ENTITY GATE_NOT IS
    PORT (A: IN STD_LOGIC; O: OUT STD_LOGIC);
END GATE_NOT;

--ARCHITECTURE DECLARATION FOR 1-BIT NOT
ARCHITECTURE Structural OF GATE_NOT IS
BEGIN
    O <= NOT A;
END Structural;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--ENTITY DECLARATION FOR 16-BIT NOT
ENTITY GATE_NOT_16 IS
	PORT (A: IN STD_LOGIC_VECTOR(15 DOWNTO 0); O: OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END GATE_NOT_16;

--ARCHITECTURE DECLARATION FOR 16-BIT NOT
ARCHITECTURE Structural OF GATE_NOT_16 IS BEGIN
	O <= NOT A;
END Structural;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--ENTITY DECLARATION FOR 1-BIT ADDER
ENTITY FULLADDER IS
	PORT (A, B, CIN: IN STD_LOGIC; O, COUT: OUT STD_LOGIC);
END FULLADDER;

--ARCHITECTURE DECLARATION FOR 1-BIT ADDER
ARCHITECTURE Structural OF FULLADDER IS
--COMPONENT THAT ARE USED NEED TO BE DECLARED AGAIN
COMPONENT GATE_XOR_3 PORT (A, B, C: IN STD_LOGIC; O: OUT STD_LOGIC);
END COMPONENT;
COMPONENT GATE_AND_2 PORT (A, B: IN STD_LOGIC; O: OUT STD_LOGIC);
END COMPONENT;
COMPONENT GATE_OR_3 PORT (A, B, C: IN STD_LOGIC; O: OUT STD_LOGIC);
END COMPONENT;
--SIGNAL TEMP STD_LOGIC
SIGNAL T1, T2, T3: STD_LOGIC;
BEGIN
	--INSTANTATE APPROPRIATE GATES
	V0: GATE_XOR_3 PORT MAP(A, B, CIN, O);
	V1: GATE_AND_2 PORT MAP(A, B, T1);
	V2: GATE_AND_2 PORT MAP(A, CIN, T2);
	V3: GATE_AND_2 PORT MAP(B, CIN, T3);
	V4: GATE_OR_3 PORT MAP(T1, T2, T3, COUT);
END Structural;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--ENTITY DECLARATION FOR 16-BIT ADDER
ENTITY FULLADDER_16 IS
	PORT (A, B: IN STD_LOGIC_VECTOR (15 DOWNTO 0); CIN: IN STD_LOGIC; O16: OUT STD_LOGIC_VECTOR (15 DOWNTO 0); V, COUT: OUT STD_LOGIC);
END FULLADDER_16;

--ARCHITECTURE DECLARATION FOR 16-BIT ADDER
ARCHITECTURE Structural OF FULLADDER_16 IS
--COMPONENTS THAT ARE USED NEED TO BE DECLARED AGAIN
COMPONENT FULLADDER PORT(A, B, CIN: IN STD_LOGIC; O, COUT: OUT STD_LOGIC);
END COMPONENT;
COMPONENT GATE_XOR PORT(A, B: IN STD_LOGIC; O: OUT STD_LOGIC);
END COMPONENT;
SIGNAL C: STD_LOGIC_VECTOR(16 DOWNTO 1);
BEGIN
	--INSTANTATE APPROPRIATE GATES & FUNCTIONS
	FA0: FULLADDER PORT MAP(A(0), B(0), CIN, O16(0), C(1));
	FA1: FULLADDER PORT MAP(A(1), B(1), C(1), O16(1), C(2));
	FA2: FULLADDER PORT MAP(A(2), B(2), C(2), O16(2), C(3));
	FA3: FULLADDER PORT MAP(A(3), B(3), C(3), O16(3), C(4));
	FA4: FULLADDER PORT MAP(A(4), B(4), C(4), O16(4), C(5));
	FA5: FULLADDER PORT MAP(A(5), B(5), C(5), O16(5), C(6));
	FA6: FULLADDER PORT MAP(A(6), B(6), C(6), O16(6), C(7));
	FA7: FULLADDER PORT MAP(A(7), B(7), C(7), O16(7), C(8));
	FA8: FULLADDER PORT MAP(A(8), B(8), C(8), O16(8), C(9));
	FA9: FULLADDER PORT MAP(A(9), B(9), C(9), O16(9), C(10));
	FA10: FULLADDER PORT MAP(A(10), B(10), C(10), O16(10), C(11));
	FA11: FULLADDER PORT MAP(A(11), B(11), C(11), O16(11), C(12));
	FA12: FULLADDER PORT MAP(A(12), B(12), C(12), O16(12), C(13));
	FA13: FULLADDER PORT MAP(A(13), B(13), C(13), O16(13), C(14));
	FA14: FULLADDER PORT MAP(A(14), B(14), C(14), O16(14), C(15));
	FA15: FULLADDER PORT MAP(A(15), B(15), C(15), O16(15), C(16));
	INST_XOR: GATE_XOR PORT MAP(C(15), C(16), V);
	--V <= C(15) XOR C(16);
	COUT <= C(16);
END Structural;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
USE ieee.numeric_std.all;

--ENTITY DECLARATION FOR 16-BIT SUBTRACTOR
ENTITY SUBTRACTOR_16 IS
	PORT(A, B: IN STD_LOGIC_VECTOR (15 DOWNTO 0); CIN: IN STD_LOGIC; O16: OUT STD_LOGIC_VECTOR (15 DOWNTO 0); V, COUT: OUT STD_LOGIC);
END SUBTRACTOR_16;

--ARCHITECTURE DECLARATION FOR 16-BIT SUBTRACTOR
ARCHITECTURE Structural OF SUBTRACTOR_16 IS
--SIGNAL TEMP STD_LOGIC_VECTOR & STD_LOGIC
SIGNAL NOT_B_RES: STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL COUT_RES: STD_LOGIC;
--COMPONENTS THAT ARE USED NEED TO BE DECLARED AGAIN
COMPONENT GATE_NOT_16 PORT (A: IN STD_LOGIC_VECTOR(15 DOWNTO 0); O: OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END COMPONENT;
COMPONENT FULLADDER_16 PORT(A, B: IN STD_LOGIC_VECTOR (15 DOWNTO 0); CIN: IN STD_LOGIC; O16: OUT STD_LOGIC_VECTOR (15 DOWNTO 0); V, COUT: OUT STD_LOGIC);
END COMPONENT;
COMPONENT GATE_NOT PORT (A: IN STD_LOGIC; O: OUT STD_LOGIC);
END COMPONENT;
BEGIN
	--INSTANTATE APPROPRIATE GATES & FUNCTIONS
	NOT_B: GATE_NOT_16 PORT MAP(B, NOT_B_RES);
	SUB: FULLADDER_16 PORT MAP(A, NOT_B_RES, CIN, O16, V, COUT_RES);
	NOT_COUT: GATE_NOT PORT MAP(COUT_RES, COUT);
END Structural;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--ENTITY DECLARATION FOR COUNTER
ENTITY COUNTER IS
	PORT(CLEAR, CLOCK : IN STD_LOGIC; Q: OUT STD_LOGIC_VECTOR(1 DOWNTO 0));
END COUNTER;

--ARCHITECTURE DECLARATION FOR COUNTER
ARCHITECTURE Structural OF COUNTER IS 
	--SIGNAL TEMP STD_LOGIC_VECTOR
	SIGNAL COUNT : STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN
	PROCESS (CLOCK)
	BEGIN
		IF (CLOCK'EVENT AND CLOCK = '1') THEN
			IF CLEAR = '1' THEN
				COUNT <= "00";
			ELSE
				COUNT <= COUNT + 1;
			END IF;
		END IF;
	END PROCESS;
	Q <= COUNT;
END Structural;

library ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

--ENTITY DECLARATION FOR 16-BIT FLIP FLOP
ENTITY REG IS
	PORT (I: IN STD_LOGIC_VECTOR(15 DOWNTO 0); EN, CLOCK: IN STD_LOGIC; O: BUFFER STD_LOGIC_VECTOR(15 DOWNTO 0));
END REG;

--ARCHITECTURE DECLARATION FOR 16-BIT FLIP FLOP
ARCHITECTURE Structural OF REG IS
BEGIN
	PROCESS (CLOCK)
	BEGIN
		IF CLOCK'EVENT AND CLOCK = '1' THEN
			IF EN = '1' THEN
				O <= I;
			END IF;
		END IF;
	END PROCESS;
END Structural;